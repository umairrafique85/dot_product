module vec_dot_product_8_treeadd_comparator (
    input logic [64-1:0] vec_a, vec_b,
    output logic [19-1:0] dot_product_bhv_treeadd_explicit, dot_product_bhv_treeadd_packed, dot_product_bhv_treadd_unpacked, vec_dot_product_8_bhv_param
);
    vec_dot_product_8_bhv_treeadd_explicit (
        .vec_a(vec_a),
        .vec_b(vec_b),
        .dot_product(dot_product_bhv_treeadd_explicit)
    );
    vec_dot_product_8_bhv_treeadd_packed (
        .vec_a(vec_a),
        .vec_b(vec_b),
        .dot_product(dot_product_bhv_treeadd_packed)
    );
    vec_dot_product_8_bhv_treeadd_unpacked (
        .vec_a(vec_a),
        .vec_b(vec_b),
        .dot_product(dot_product_bhv_treeadd_unpacked)
    );
    vector_dot_product_8_bhv_treeadd_param (
        .vec_a(vec_a),
        .vec_b(vec_b),
        .dot_product(dot_product_bhv_treeadd_param)
    );
endmodule

// Claude
// Using explicit tree-based adder
module vec_dot_product_8_bhv_treeadd_explicit (
    input  logic [64-1:0] vec_a, vec_b,
    output logic [19-1:0] dot_product
);
    // Break vectors into individual bytes for clarity
    logic [7:0] a_bytes [7:0];
    logic [7:0] b_bytes [7:0];
    logic [15:0] products [7:0];

    // Extract bytes explicitly
    genvar i;
    generate
        for (i = 0; i < 8; i++) begin : proc_extract_multiply
            assign a_bytes[i] = vec_a[i*8 +: 8];
            assign b_bytes[i] = vec_b[i*8 +: 8];
            assign products[i] = a_bytes[i] * b_bytes[i];
        end
    endgenerate

    // Tree-based addition for better timing
    logic [16:0] sum_level1 [3:0];
    logic [17:0] sum_level2 [1:0];

    assign sum_level1[0] = products[0] + products[1];
    assign sum_level1[1] = products[2] + products[3];
    assign sum_level1[2] = products[4] + products[5];
    assign sum_level1[3] = products[6] + products[7];

    assign sum_level2[0] = sum_level1[0] + sum_level1[1];
    assign sum_level2[1] = sum_level1[2] + sum_level1[3];

    assign dot_product = sum_level2[0] + sum_level2[1];
endmodule

// Same target, generate block, packed intermediary vectors
module vec_dot_product_8_bhv_treeadd_packed (
    input logic [64-1:0] vec_a, vec_b,
    output [19-1:0] dot_product
);

    logic [15:0] products [8-1:0]; // Array of products

    genvar i;
    generate
        for (i = 0; i < 8; i++) begin: proc_multiply
            assign products[i] = vec_a[i*8 +: 8] * vec_b[i*8 +: 8];
        end
    endgenerate

    logic [17*4-1:0] sum_level1;
    logic [18*2-1:0] sum_level2;

    genvar j;
    generate
        for (j = 0; j < 4; j++) begin: proc_add_stage_1
            assign sum_level1[j*17 +: 17] = products[j*2] + products[j*2+1];
        end
    endgenerate

    genvar k;
    generate
        for (k = 0; k < 2; k++) begin: proc_add_state_2
            assign sum_level2[k*18 +: 18] = sum_level1[k*2*17 +: 17] + sum_level1[(k*2+1)*17 +: 17];
        end
    endgenerate

    assign dot_product = sum_level2[36-1:18] + sum_level2[18-1:0];
endmodule

// Generate blocks for intermediary addition steps, unpacked arrays
module vec_dot_product_8_bhv_treeadd_unpacked (
    input  logic [63:0] vec_a, vec_b, // can use packed 2D here as well
    output logic [18:0] dot_product
);
    logic [15:0] products [8];
    logic [16:0] sum_l1 [4];
    logic [17:0] sum_l2 [2];

    genvar i, j, k;
    generate
        for (i = 0; i < 8; i++) begin : gen_mult
            assign products[i] = vec_a[i*8 +: 8] * vec_b[i*8 +: 8]; // if using packed 2D, just use [i]
        end

        for (j = 0; j < 4; j++) begin : gen_l1
            assign sum_l1[j] = products[2*j] + products[2*j+1];
        end

        for (k = 0; k < 2; k++) begin : gen_l2
            assign sum_l2[k] = sum_l1[2*k] + sum_l1[2*k+1];
        end
    endgenerate

    assign dot_product = sum_l2[0] + sum_l2[1];
endmodule

// Claude: PARAMETERIZED VERSION: Most flexible and reusable
// using function for treeadder
// ############## DOES NOT CREATE TREEADDER LIKE CLAUDE CLAIMED ###############
module vector_dot_product_8_bhv_treeadd_param #(
    parameter int NUM_ELEMENTS = 8,
    parameter int ELEMENT_WIDTH = 8,
    parameter int VECTOR_WIDTH = NUM_ELEMENTS * ELEMENT_WIDTH
) (
    input  logic [ELEMENT_WIDTH-1:0][NUM_ELEMENTS-1:0] vec_a, vec_b,
    output logic [$clog2(NUM_ELEMENTS * (2**ELEMENT_WIDTH)**2)-1:0] dot_product
);
    // Calculate product width: element_width * 2
    localparam int PRODUCT_WIDTH = ELEMENT_WIDTH * 2;

    logic [ELEMENT_WIDTH-1:0] a_elements [NUM_ELEMENTS-1:0];
    logic [ELEMENT_WIDTH-1:0] b_elements [NUM_ELEMENTS-1:0];
    logic [PRODUCT_WIDTH-1:0] products [NUM_ELEMENTS-1:0];

    // Extract elements and compute products
    genvar i;
    generate
        for (i = 0; i < NUM_ELEMENTS; i++) begin : gen_dot_product
            assign products[i] = vec_a[i] * vec_b[i];
        end
    endgenerate

    // Recursive tree summation function
    function automatic logic [$clog2(NUM_ELEMENTS * (2**ELEMENT_WIDTH)**2)-1:0] sum_products;
        input logic [PRODUCT_WIDTH-1:0] prods [NUM_ELEMENTS-1:0];
        logic [$clog2(NUM_ELEMENTS * (2**ELEMENT_WIDTH)**2)-1:0] result;
        begin
            result = 0;
            for (int j = 0; j < NUM_ELEMENTS; j++) begin
                result = result + prods[j];
            end
            sum_products = result;
        end
    endfunction

    assign dot_product = sum_products(products);
endmodule

// Claude: Using systemverilog array sum function
// ################# Not compiling. Apparently needs IP########################
module vec_dot_product_8_bhv_funadd (
    input  logic [8-1:0][8-1:0] vec_a, vec_b,  // 2D packed array
    output logic [19-1:0]     dot_product
);
    // Using SystemVerilog reduction
    logic [15:0] products [8];

    always_comb begin
        for (int i = 0; i < 8; i++) begin
            products[i] = vec_a[i] * vec_b[i];
        end

        // Could use array reduction functions
        dot_product = products.sum();  // SystemVerilog array method
    end
endmodule
